`timescale 1ns / 1ps 

module top(
           input  sw,
           output led
           );
   assign led = sw;
endmodule
